module singlecycle(
    input resetl,
    input [63:0] startpc,
    output reg [63:0] currentpc,
    output [63:0] dmemout,
    input CLK
);

    // Next PC connections
    wire [63:0] nextpc;       // The next PC, to be updated on clock cycle

    // Instruction Memory connections
    wire [31:0] instruction;  // The current instruction

    // Parts of instruction
    wire [4:0] rd;            // The destination register
    wire [4:0] rm;            // Operand 1
    wire [4:0] rn;            // Operand 2
    wire [10:0] opcode;
   

    // Control wires
    wire reg2loc;
    wire alusrc;
    wire mem2reg;
    wire regwrite;
    wire memread;
    wire memwrite;
    wire branch;
    wire uncond_branch;
    wire [3:0] aluctrl;
    wire        move;
    wire [2:0] signop;

    // Register file connections
    wire [63:0] regoutA;     // Output A
    wire [63:0] regoutB;     // Output B
   wire [63:0] 	writedata;   //2x1 move mux input
   wire [63:0] 	finalwrite;  //Write data input
   

    // ALU connections
   wire [63:0] 	b_input;    //Defining the b_input between mux and ALU
    wire [63:0] aluout;
    wire zero;

    // Sign Extender connections
   wire [25:0] signext;    //Defining input for sign extend module
    wire [63:0] extimm;    //Sign extender output

    // PC update logic
    always @(negedge CLK)
    begin
        if (resetl)
            currentpc <= nextpc;
        else
            currentpc <= startpc;
    end

    // Parts of instruction
    assign rd = instruction[4:0];
    assign rm = instruction[9:5];
    assign rn = reg2loc ? instruction[4:0] : instruction[20:16];  //Mux before Read register 2
    assign opcode = instruction[31:21];
   assign signext = instruction[25:0];     //Setting signext to be first 26 bits of instruction
   
   

    InstructionMemory imem(
			   .Data(instruction),
			   .Address(currentpc)
    );

    control control(
		    .reg2loc(reg2loc),
		    .alusrc(alusrc),
		    .mem2reg(mem2reg),
		    .regwrite(regwrite),
		    .memread(memread),
		    .memwrite(memwrite),
		    .branch(branch),
		    .uncond_branch(uncond_branch),
		    .move(move),
		    .aluop(aluctrl),
		    .signop(signop),
		    .opcode(opcode)
    );

    /*
    * Connect the remaining datapath elements below.
    * Do not forget any additional multiplexers that may be required.
    */
   RegisterFile RegisterFile(
			     .BusA(regoutA),
			     .BusB(regoutB),
			     .BusW(finalwrite),
			     .RA(rm),
			     .RB(rn),
			     .RW(rd),
			     .RegWr(regwrite),
			     .Clk(CLK)   
			     );

   SignExtender SignExtender(
			     .BusImm(extimm),
			     .Imm26(signext),
			     .Ctrl(signop)
			     );
   	     
   assign b_input = alusrc ? extimm : regoutB;    //MUX taking Read data 2 and Sign Extended value as inputs, output is an input to the ALU.
   assign finalwrite = move ? extimm : writedata; //Mux that writes sign extended MOVZ if move is true.
   
   ALU ALU(
	   .BusW(aluout),
	   .BusA(regoutA),
	   .BusB(b_input),
	   .ALUCtrl(aluctrl),
	   .Zero(zero)
	   );

   NextPClogic NextPClogic(
		      .NextPC(nextpc),
		      .CurrentPC(currentpc),
		      .SignExtImm64(extimm),
		      .Branch(branch),
		      .ALUZero(zero),
		      .Uncondbranch(uncond_branch)
		      );

   DataMemory DataMemory(
			 .ReadData(dmemout),
			 .Address(aluout),
			 .WriteData(regoutB),
			 .MemoryRead(memread),
			 .MemoryWrite(memwrite),
			 .Clock(CLK)
			 );
   
   assign writedata = mem2reg ? dmemout : aluout;  //Mux that takes read data and aluout as inputs, output is the input to write data in register file.
   
   
endmodule

